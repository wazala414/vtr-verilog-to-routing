//A simple cricuit which blinks an LED on and off periodically
module null_arch(output o);
    wire a;
    //o <= null;
endmodule
